`default_nettype wire
`include "mycpu.h"

module id_stage(
    input                          clk           ,
    input                          reset         ,
    //allowin
    input                          es_allowin    ,
    output                         ds_allowin    ,
    //from fs
    input                          fs_to_ds_valid,
    input  [`FS_TO_DS_BUS_WD -1:0] fs_to_ds_bus  ,
    //to es
    output                         ds_to_es_valid,
    output [`DS_TO_ES_BUS_WD -1:0] ds_to_es_bus  ,
    //to fs
    output [`BR_BUS_WD       -1:0] br_bus        ,
    //to rf: for write back
    input  [`WS_TO_RF_BUS_WD -1:0] ws_to_rf_bus,
    //receive later stages' forward dest
    input [4:0] es_fwd_dest,
    input [4:0] ms_fwd_dest,
    input [4:0] ws_fwd_dest,
    //reveive later stages' forward result
    input [31:0] es_fwd_res,
    input [31:0] ms_fwd_res,
    input [31:0] ws_fwd_res,
    input       es_ld
);

reg         ds_valid   ;
wire        ds_ready_go;

reg  [`FS_TO_DS_BUS_WD -1:0] fs_to_ds_bus_r;

wire [31:0] ds_inst;
wire [31:0] ds_pc  ;
assign {ds_inst,
        ds_pc  } = fs_to_ds_bus_r;

wire        rf_we   ;
wire [ 4:0] rf_waddr;
wire [31:0] rf_wdata;
assign {rf_we   ,  //37:37
        rf_waddr,  //36:32
        rf_wdata   //31:0
       } = ws_to_rf_bus;

wire        br_taken;
wire [31:0] br_target;

wire        ld_signed;
wire        ls_width_h;
wire        ls_width_b;
wire        op_need_div;
wire        op_need_mul;
wire        md_signed;
wire        md_high;
wire [11:0] alu_op;
wire        load_op;
wire        src1_is_pc;
wire        src2_is_imm;
wire        dst_is_r1;
wire        gr_we;
wire        mem_we;
wire        src_reg_is_rd;
wire [4: 0] dest;
wire [31:0] rj_value;
wire [31:0] rkd_value;
wire [31:0] ds_imm;
wire [31:0] br_offs;
wire [31:0] jirl_offs;

wire [ 5:0] op_31_26;
wire [ 3:0] op_25_22;
wire [ 1:0] op_21_20;
wire [ 4:0] op_19_15;
wire [ 4:0] rd;
wire [ 4:0] rj;
wire [ 4:0] rk;
wire [11:0] i12;
wire [19:0] i20;
wire [15:0] i16;
wire [25:0] i26;

wire [63:0] op_31_26_d;
wire [15:0] op_25_22_d;
wire [ 3:0] op_21_20_d;
wire [31:0] op_19_15_d;

wire        inst_add_w;
wire        inst_sub_w;
wire        inst_slt;
wire        inst_sltu;
wire        inst_nor;
wire        inst_and;
wire        inst_or;
wire        inst_xor;
wire        inst_slli_w;
wire        inst_srli_w;
wire        inst_srai_w;
wire        inst_addi_w;
wire        inst_ld_w;
wire        inst_st_w;
wire        inst_jirl;
wire        inst_b;
wire        inst_bl;
wire        inst_beq;
wire        inst_bne;
wire        inst_lu12i_w;
//new
wire        inst_slti;
wire        inst_sltui;
wire        inst_andi;
wire        inst_ori;
wire        inst_xori;
wire        inst_sll;
wire        inst_srl;
wire        inst_sra;
wire        in_pcaddu12i;
// mul div
wire        inst_mul_w;
wire        inst_mulh_w;
wire        inst_mulh_wu;
wire        inst_div_w;
wire        inst_mod_w;
wire        inst_div_wu;
wire        inst_mod_wu;
//new exp11 branch
wire        inst_blt;
wire        inst_bge;
wire        inst_bltu;
wire        inst_bgeu;
wire        inst_is_branch;  //branch inst set
//new exp11 load store
wire        inst_ld_b;
wire        inst_ld_h;
wire        inst_ld_bu;
wire        inst_ld_hu;
wire        inst_st_b;
wire        inst_st_h;

wire        need_ui5;
wire        need_ui12;  //new
wire        need_si12;
wire        need_si16;
wire        need_si20;
wire        need_si26;
wire        src2_is_4;

wire [ 4:0] rf_raddr1;
wire [31:0] rf_rdata1;
wire [ 4:0] rf_raddr2;
wire [31:0] rf_rdata2;

wire        rj_eq_rd;
wire        rj_lt_rd;
wire        rj_lt_ud;

assign ld_signed    = inst_ld_b | inst_ld_h ;
assign ls_width_h   = inst_st_h | inst_ld_h | inst_ld_hu;
assign ls_width_b   = inst_st_b | inst_ld_b | inst_ld_bu;
assign load_op      = inst_ld_w | inst_ld_b | inst_ld_h | inst_ld_bu | inst_ld_hu;
assign mem_we       = inst_st_w | inst_st_h | inst_st_b ;
assign gr_we        = ~mem_we & ~inst_is_branch & ~inst_b;
assign dst_is_r1    = inst_bl;
assign dest         = dst_is_r1 ? 5'd1 : rd;

assign ds_to_es_bus = {ld_signed   ,  //156:156
                       ls_width_h  ,  //155:155
                       ls_width_b  ,  //154:154
                       op_need_div ,  //153:153
                       op_need_mul ,  //152:152
                       md_signed   ,  //151:151
                       md_high     ,  //150:150
                       alu_op      ,  //149:138
                       load_op     ,  //137:137
                       src1_is_pc  ,  //136:136
                       src2_is_imm ,  //135:135
                       gr_we       ,  //134:134
                       mem_we      ,  //133:133
                       dest        ,  //132:128
                       ds_imm      ,  //127:96
                       rj_value    ,  //95 :64
                       rkd_value   ,  //63 :32
                       ds_pc          //31 :0
                      };

wire rj_comparable;
wire rk_comparable;
wire rd_comparable;
wire rj_conflict;
wire rk_conflict;
wire rd_conflict;
wire es_ld_wait;

assign rj_comparable = (rj!=5'd0) && ~(need_si20 | need_si26);
assign rk_comparable = (rk!=5'd0) && ~(src2_is_imm | inst_b | inst_is_branch);
assign rd_comparable = (rd!=5'd0) && src_reg_is_rd;
assign rj_conflict = rj_comparable && rj == es_fwd_dest;
assign rk_conflict = rk_comparable && rk == es_fwd_dest;
assign rd_conflict = rd_comparable && rd == es_fwd_dest;
assign es_ld_wait = (rj_conflict || rk_conflict || rd_conflict) && es_ld;

assign ds_ready_go    = ~es_ld_wait;
assign ds_allowin     = !ds_valid || ds_ready_go && es_allowin;
assign ds_to_es_valid = ds_valid && ds_ready_go;
always @(posedge clk) begin
    if (reset) begin
        ds_valid <= 1'b0;
    end
    else if (br_taken) begin
        ds_valid <= 1'b0;
    end
    else if (es_allowin) begin
        ds_valid <= fs_to_ds_valid;
    end
    if (fs_to_ds_valid && ds_allowin) begin
        fs_to_ds_bus_r <= fs_to_ds_bus;
    end
end

assign op_31_26  = ds_inst[31:26];
assign op_25_22  = ds_inst[25:22];
assign op_21_20  = ds_inst[21:20];
assign op_19_15  = ds_inst[19:15];

assign rd   = ds_inst[ 4: 0];
assign rj   = ds_inst[ 9: 5];
assign rk   = ds_inst[14:10];

assign i12  = ds_inst[21:10];
assign i20  = ds_inst[24: 5];
assign i16  = ds_inst[25:10];
assign i26  = {ds_inst[ 9: 0], ds_inst[25:10]};

decoder #(.WIDTH(6)) u_dec6(.in(op_31_26), .out(op_31_26_d));
decoder #(.WIDTH(4)) u_dec4(.in(op_25_22), .out(op_25_22_d));
decoder #(.WIDTH(2)) u_dec2(.in(op_21_20), .out(op_21_20_d));
decoder #(.WIDTH(5)) u_dec5(.in(op_19_15), .out(op_19_15_d));

assign inst_add_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h00];
assign inst_sub_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h02];
assign inst_slt    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h04];
assign inst_sltu   = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h05];
assign inst_nor    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h08];
assign inst_and    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h09];
assign inst_or     = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0a];
assign inst_xor    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0b];
assign inst_slli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h01];
assign inst_srli_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h09];
assign inst_srai_w = op_31_26_d[6'h00] & op_25_22_d[4'h1] & op_21_20_d[2'h0] & op_19_15_d[5'h11];
assign inst_addi_w = op_31_26_d[6'h00] & op_25_22_d[4'ha];
assign inst_ld_w   = op_31_26_d[6'h0a] & op_25_22_d[4'h2];
assign inst_st_w   = op_31_26_d[6'h0a] & op_25_22_d[4'h6];
assign inst_jirl   = op_31_26_d[6'h13];
assign inst_b      = op_31_26_d[6'h14];
assign inst_bl     = op_31_26_d[6'h15];
assign inst_beq    = op_31_26_d[6'h16];
assign inst_bne    = op_31_26_d[6'h17];
assign inst_lu12i_w= op_31_26_d[6'h05] & ~ds_inst[25];
//new inst
assign inst_slti   = op_31_26_d[6'h00] & op_25_22_d[4'h8];
assign inst_sltui  = op_31_26_d[6'h00] & op_25_22_d[4'h9];
assign inst_andi   = op_31_26_d[6'h00] & op_25_22_d[4'hd];
assign inst_ori    = op_31_26_d[6'h00] & op_25_22_d[4'he];
assign inst_xori   = op_31_26_d[6'h00] & op_25_22_d[4'hf];
assign inst_sll    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0e];
assign inst_srl    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h0f];
assign inst_sra    = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h10];
assign in_pcaddu12i= op_31_26_d[6'h07] & ~ds_inst[25];
//mul, div
assign inst_mul_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h18];
assign inst_mulh_w = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h19];
assign inst_mulh_wu= op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h1] & op_19_15_d[5'h1a];
assign inst_div_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h00];
assign inst_mod_w  = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h01];
assign inst_div_wu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h02];
assign inst_mod_wu = op_31_26_d[6'h00] & op_25_22_d[4'h0] & op_21_20_d[2'h2] & op_19_15_d[5'h03];
// new exp11 branch
assign inst_blt    = op_31_26_d[6'h18];
assign inst_bge    = op_31_26_d[6'h19];
assign inst_bltu   = op_31_26_d[6'h1a];
assign inst_bgeu   = op_31_26_d[6'h1b];
// new exp11 load store
assign inst_ld_b   = op_31_26_d[6'h0a] & op_25_22_d[4'h0];
assign inst_ld_h   = op_31_26_d[6'h0a] & op_25_22_d[4'h1];
assign inst_ld_bu  = op_31_26_d[6'h0a] & op_25_22_d[4'h8];
assign inst_ld_hu  = op_31_26_d[6'h0a] & op_25_22_d[4'h9];
assign inst_st_b   = op_31_26_d[6'h0a] & op_25_22_d[4'h4];
assign inst_st_h   = op_31_26_d[6'h0a] & op_25_22_d[4'h5];

assign inst_is_branch = inst_beq  | inst_bne  | inst_blt   | inst_bge  | inst_bltu | inst_bgeu;

assign alu_op[ 0] = inst_add_w | inst_addi_w | load_op | mem_we
                  | inst_jirl | inst_bl | in_pcaddu12i;
assign alu_op[ 1] = inst_sub_w;
assign alu_op[ 2] = inst_slt | inst_slti;
assign alu_op[ 3] = inst_sltu | inst_sltui;
assign alu_op[ 4] = inst_and | inst_andi;
assign alu_op[ 5] = inst_nor;
assign alu_op[ 6] = inst_or | inst_ori;
assign alu_op[ 7] = inst_xor | inst_xori;
assign alu_op[ 8] = inst_slli_w | inst_sll;
assign alu_op[ 9] = inst_srli_w | inst_srl;
assign alu_op[10] = inst_srai_w | inst_sra;
assign alu_op[11] = inst_lu12i_w;

assign op_need_mul= inst_mul_w | inst_mulh_w  | inst_mulh_wu;
assign op_need_div= inst_div_w | inst_div_wu  | inst_mod_w  | inst_mod_wu;
assign md_signed  = inst_mulh_w| inst_div_w   | inst_mod_w  ;
assign md_high    = inst_mulh_w| inst_mulh_wu | inst_div_w  | inst_div_wu;

assign need_ui5   = inst_slli_w | inst_srli_w | inst_srai_w;
assign need_ui12  = inst_andi   | inst_ori    | inst_xori;
assign need_si12  = inst_addi_w | load_op     | mem_we      | inst_sltui | inst_slti;
assign need_si16  = inst_jirl   | inst_is_branch;
assign need_si20  = inst_lu12i_w| in_pcaddu12i;
assign need_si26  = inst_b      | inst_bl;
assign src2_is_4  = inst_jirl   | inst_bl;

//TODO: rectify
assign ds_imm = src2_is_4 ? 32'h4                      :
                need_si20 ? {i20[19:0]    ,     12'b0} :
                need_si12 ? {{20{i12[11]}}, i12[11:0]} :
  /*need_ui5 || need_ui12 */{20'b0        , i12[11:0]} ;

assign br_offs = need_si26 ? {{ 4{i26[25]}}, i26[25:0], 2'b0} :
               /*need_si16*/ {{14{i16[15]}}, i16[15:0], 2'b0} ;

assign jirl_offs = {{14{i16[15]}}, i16[15:0], 2'b0};

assign src_reg_is_rd = inst_is_branch | mem_we;

assign src1_is_pc    = inst_jirl | inst_bl | in_pcaddu12i;

assign src2_is_imm   = inst_slli_w |
                       inst_srli_w |
                       inst_srai_w |
                       inst_addi_w |
                       load_op     |
                       mem_we      |
                       inst_lu12i_w|
                       inst_jirl   |
                       inst_bl     |
                       inst_slti   |
                       inst_sltui  |
                       inst_ori    |
                       inst_andi   |
                       inst_xori   |
                       in_pcaddu12i;


assign rf_raddr1 = rj;
assign rf_raddr2 = src_reg_is_rd ? rd :rk;
regfile u_regfile(
    .clk    (clk      ),
    .raddr1 (rf_raddr1),
    .rdata1 (rf_rdata1),
    .raddr2 (rf_raddr2),
    .rdata2 (rf_rdata2),
    .we     (rf_we    ),
    .waddr  (rf_waddr ),
    .wdata  (rf_wdata )
    );


assign rj_value  = rj_comparable ? 
                  (rj == es_fwd_dest) ? es_fwd_res :
                  (rj == ms_fwd_dest) ? ms_fwd_res :
                  (rj == ws_fwd_dest) ? ws_fwd_res : rf_rdata1
                  : rf_rdata1;
assign rkd_value = (rd_comparable || rk_comparable) ?
                   (rf_raddr2 == es_fwd_dest) ? es_fwd_res :
                   (rf_raddr2 == ms_fwd_dest) ? ms_fwd_res :
                   (rf_raddr2 == ws_fwd_dest) ? ws_fwd_res : rf_rdata2
                  : rf_rdata2;

assign rj_eq_rd = (rj_value == rkd_value);
assign rj_lt_ud = (rj_value <  rkd_value);
assign rj_lt_rd = ($signed(rj_value) < $signed(rkd_value));

assign br_taken = (   inst_beq  &&  rj_eq_rd  && ds_ready_go
                   || inst_bne  && !rj_eq_rd  && ds_ready_go
                   || inst_blt  &&  rj_lt_rd  && ds_ready_go
                   || inst_bltu &&  rj_lt_ud  && ds_ready_go
                   || inst_bge  && !rj_lt_rd  && ds_ready_go
                   || inst_bgeu && !rj_lt_ud  && ds_ready_go
                   || inst_jirl
                   || inst_bl
                   || inst_b
                  ) && ds_valid;

assign br_target = (inst_is_branch|| inst_bl || inst_b) ? (ds_pc + br_offs)
                                         /*inst_jirl*/  : (rj_value + jirl_offs);

assign br_bus       ={br_taken  , br_target};

endmodule
